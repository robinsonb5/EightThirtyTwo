
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.rom_pkg.all;

entity dhry_1_rom is
generic
	(
		maxAddrBitBRAM : natural := maxAddrBitBRAMLimit;
		BYTE_WIDTH : natural := 8;
		BYTES : natural := 4
--		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_soc : in toROM;
	to_soc : out fromROM
);
end entity;

architecture rtl of dhry_1_rom is

	alias be1 is from_soc.memAByteSel;
	alias we1 is from_soc.memAWriteEnable;
	alias data_in1 is from_soc.memAWrite;
	signal addr1 : integer range 0 to 2**maxAddrBitBRAM-1;
	alias data_out1 is to_soc.memARead;

	--  build up 2D array to hold the memory
	type word_t is array (0 to BYTES-1) of std_logic_vector(BYTE_WIDTH-1 downto 0);
	type ram_t is array (0 to 2 ** (maxAddrBitBRAM-1) - 1) of word_t;

	signal ram : ram_t:=
	(
     0 => (x"04",x"87",x"c9",x"01"),
     1 => (x"cf",x"03",x"87",x"cc"),
     2 => (x"87",x"fd",x"00",x"87"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"36",x"27",x"4f",x"00"),
     5 => (x"4f",x"00",x"00",x"00"),
     6 => (x"0e",x"1e",x"18",x"0e"),
     7 => (x"00",x"00",x"44",x"27"),
     8 => (x"48",x"26",x"0f",x"00"),
     9 => (x"08",x"26",x"80",x"ff"),
    10 => (x"c0",x"e0",x"c0",x"4f"),
    11 => (x"02",x"e9",x"27",x"4e"),
    12 => (x"00",x"0f",x"00",x"00"),
    13 => (x"d0",x"c0",x"87",x"fd"),
    14 => (x"43",x"27",x"4e",x"c0"),
    15 => (x"0f",x"00",x"00",x"00"),
    16 => (x"4f",x"87",x"fd",x"00"),
    17 => (x"0e",x"1e",x"18",x"0e"),
    18 => (x"80",x"ff",x"48",x"26"),
    19 => (x"1e",x"4f",x"08",x"26"),
    20 => (x"ff",x"1e",x"1e",x"72"),
    21 => (x"48",x"6a",x"4a",x"c0"),
    22 => (x"c4",x"98",x"c0",x"c4"),
    23 => (x"02",x"6e",x"58",x"a6"),
    24 => (x"cc",x"87",x"f3",x"ff"),
    25 => (x"66",x"cc",x"7a",x"66"),
    26 => (x"4a",x"26",x"26",x"48"),
    27 => (x"5e",x"0e",x"4f",x"26"),
    28 => (x"5d",x"5c",x"5b",x"5a"),
    29 => (x"4d",x"66",x"d4",x"0e"),
    30 => (x"4b",x"15",x"4c",x"c0"),
    31 => (x"c0",x"02",x"9b",x"73"),
    32 => (x"4a",x"73",x"87",x"d6"),
    33 => (x"4f",x"27",x"1e",x"72"),
    34 => (x"0f",x"00",x"00",x"00"),
    35 => (x"84",x"c1",x"86",x"c4"),
    36 => (x"9b",x"73",x"4b",x"15"),
    37 => (x"87",x"ea",x"ff",x"05"),
    38 => (x"4d",x"26",x"48",x"74"),
    39 => (x"4b",x"26",x"4c",x"26"),
    40 => (x"4f",x"26",x"4a",x"26"),
    41 => (x"5b",x"5a",x"5e",x"0e"),
    42 => (x"1e",x"0e",x"5d",x"5c"),
    43 => (x"27",x"4d",x"66",x"d8"),
    44 => (x"00",x"00",x"16",x"30"),
    45 => (x"27",x"49",x"76",x"4b"),
    46 => (x"00",x"00",x"0e",x"70"),
    47 => (x"75",x"4c",x"c0",x"79"),
    48 => (x"a9",x"b7",x"c0",x"49"),
    49 => (x"87",x"ce",x"c0",x"03"),
    50 => (x"27",x"1e",x"ed",x"c0"),
    51 => (x"00",x"00",x"00",x"4f"),
    52 => (x"c0",x"86",x"c4",x"0f"),
    53 => (x"9d",x"75",x"8d",x"0d"),
    54 => (x"87",x"c6",x"c0",x"05"),
    55 => (x"c0",x"53",x"f0",x"c0"),
    56 => (x"9d",x"75",x"87",x"f6"),
    57 => (x"87",x"f0",x"c0",x"02"),
    58 => (x"1e",x"72",x"49",x"75"),
    59 => (x"4a",x"66",x"e4",x"c0"),
    60 => (x"00",x"0b",x"f0",x"27"),
    61 => (x"4a",x"26",x"0f",x"00"),
    62 => (x"4a",x"72",x"4a",x"71"),
    63 => (x"53",x"12",x"82",x"6e"),
    64 => (x"1e",x"72",x"49",x"75"),
    65 => (x"4a",x"66",x"e4",x"c0"),
    66 => (x"00",x"0b",x"f0",x"27"),
    67 => (x"4a",x"26",x"0f",x"00"),
    68 => (x"9d",x"75",x"4d",x"70"),
    69 => (x"87",x"d0",x"ff",x"05"),
    70 => (x"30",x"27",x"49",x"73"),
    71 => (x"b7",x"00",x"00",x"16"),
    72 => (x"e1",x"c0",x"02",x"a9"),
    73 => (x"dc",x"8b",x"c1",x"87"),
    74 => (x"97",x"49",x"bf",x"a6"),
    75 => (x"66",x"dc",x"51",x"6b"),
    76 => (x"c0",x"80",x"c1",x"48"),
    77 => (x"c1",x"58",x"a6",x"e0"),
    78 => (x"27",x"49",x"73",x"84"),
    79 => (x"00",x"00",x"16",x"30"),
    80 => (x"ff",x"05",x"a9",x"b7"),
    81 => (x"a6",x"dc",x"87",x"df"),
    82 => (x"51",x"c0",x"49",x"bf"),
    83 => (x"26",x"26",x"48",x"74"),
    84 => (x"26",x"4c",x"26",x"4d"),
    85 => (x"26",x"4a",x"26",x"4b"),
    86 => (x"5a",x"5e",x"0e",x"4f"),
    87 => (x"0e",x"5d",x"5c",x"5b"),
    88 => (x"76",x"4c",x"c0",x"1e"),
    89 => (x"dc",x"79",x"c0",x"49"),
    90 => (x"66",x"d8",x"4b",x"a6"),
    91 => (x"48",x"66",x"d8",x"4a"),
    92 => (x"a6",x"dc",x"80",x"c1"),
    93 => (x"d8",x"4d",x"12",x"58"),
    94 => (x"75",x"2d",x"b7",x"35"),
    95 => (x"d7",x"c4",x"02",x"9d"),
    96 => (x"c3",x"02",x"6e",x"87"),
    97 => (x"49",x"76",x"87",x"e1"),
    98 => (x"4a",x"75",x"79",x"c0"),
    99 => (x"e3",x"c1",x"49",x"75"),
   100 => (x"e5",x"c2",x"02",x"a9"),
   101 => (x"c1",x"49",x"72",x"87"),
   102 => (x"c0",x"02",x"a9",x"e4"),
   103 => (x"49",x"72",x"87",x"de"),
   104 => (x"02",x"a9",x"ec",x"c1"),
   105 => (x"72",x"87",x"cc",x"c2"),
   106 => (x"a9",x"f3",x"c1",x"49"),
   107 => (x"87",x"ea",x"c1",x"02"),
   108 => (x"f8",x"c1",x"49",x"72"),
   109 => (x"f2",x"c0",x"02",x"a9"),
   110 => (x"87",x"d3",x"c2",x"87"),
   111 => (x"80",x"27",x"1e",x"ca"),
   112 => (x"1e",x"00",x"00",x"16"),
   113 => (x"4a",x"73",x"83",x"c4"),
   114 => (x"1e",x"6a",x"8a",x"c4"),
   115 => (x"00",x"00",x"a4",x"27"),
   116 => (x"86",x"cc",x"0f",x"00"),
   117 => (x"4c",x"74",x"4a",x"70"),
   118 => (x"80",x"27",x"84",x"72"),
   119 => (x"1e",x"00",x"00",x"16"),
   120 => (x"00",x"00",x"6e",x"27"),
   121 => (x"86",x"c4",x"0f",x"00"),
   122 => (x"d0",x"87",x"d6",x"c2"),
   123 => (x"16",x"80",x"27",x"1e"),
   124 => (x"c4",x"1e",x"00",x"00"),
   125 => (x"c4",x"4a",x"73",x"83"),
   126 => (x"27",x"1e",x"6a",x"8a"),
   127 => (x"00",x"00",x"00",x"a4"),
   128 => (x"70",x"86",x"cc",x"0f"),
   129 => (x"72",x"4c",x"74",x"4a"),
   130 => (x"16",x"80",x"27",x"84"),
   131 => (x"27",x"1e",x"00",x"00"),
   132 => (x"00",x"00",x"00",x"6e"),
   133 => (x"c1",x"86",x"c4",x"0f"),
   134 => (x"83",x"c4",x"87",x"e7"),
   135 => (x"8a",x"c4",x"4a",x"73"),
   136 => (x"6e",x"27",x"1e",x"6a"),
   137 => (x"0f",x"00",x"00",x"00"),
   138 => (x"4a",x"70",x"86",x"c4"),
   139 => (x"84",x"72",x"4c",x"74"),
   140 => (x"76",x"87",x"ce",x"c1"),
   141 => (x"c1",x"79",x"c1",x"49"),
   142 => (x"83",x"c4",x"87",x"c7"),
   143 => (x"8a",x"c4",x"4a",x"73"),
   144 => (x"4f",x"27",x"1e",x"6a"),
   145 => (x"0f",x"00",x"00",x"00"),
   146 => (x"84",x"c1",x"86",x"c4"),
   147 => (x"c0",x"87",x"f2",x"c0"),
   148 => (x"4f",x"27",x"1e",x"e5"),
   149 => (x"0f",x"00",x"00",x"00"),
   150 => (x"1e",x"75",x"86",x"c4"),
   151 => (x"00",x"00",x"4f",x"27"),
   152 => (x"86",x"c4",x"0f",x"00"),
   153 => (x"75",x"87",x"da",x"c0"),
   154 => (x"a9",x"e5",x"c0",x"49"),
   155 => (x"87",x"c7",x"c0",x"05"),
   156 => (x"79",x"c1",x"49",x"76"),
   157 => (x"75",x"87",x"ca",x"c0"),
   158 => (x"00",x"4f",x"27",x"1e"),
   159 => (x"c4",x"0f",x"00",x"00"),
   160 => (x"4a",x"66",x"d8",x"86"),
   161 => (x"c1",x"48",x"66",x"d8"),
   162 => (x"58",x"a6",x"dc",x"80"),
   163 => (x"35",x"d8",x"4d",x"12"),
   164 => (x"9d",x"75",x"2d",x"b7"),
   165 => (x"87",x"e9",x"fb",x"05"),
   166 => (x"26",x"26",x"48",x"74"),
   167 => (x"26",x"4c",x"26",x"4d"),
   168 => (x"26",x"4a",x"26",x"4b"),
   169 => (x"5a",x"5e",x"0e",x"4f"),
   170 => (x"ff",x"0e",x"5c",x"5b"),
   171 => (x"4b",x"68",x"48",x"c8"),
   172 => (x"b7",x"d8",x"4a",x"73"),
   173 => (x"9a",x"ff",x"c3",x"2a"),
   174 => (x"b7",x"c8",x"4c",x"73"),
   175 => (x"c0",x"fc",x"cf",x"2c"),
   176 => (x"74",x"4a",x"72",x"9c"),
   177 => (x"c8",x"4c",x"73",x"b2"),
   178 => (x"f0",x"ff",x"c0",x"34"),
   179 => (x"72",x"9c",x"c0",x"c0"),
   180 => (x"d8",x"b2",x"74",x"4a"),
   181 => (x"c0",x"fc",x"cf",x"33"),
   182 => (x"72",x"9b",x"c0",x"c0"),
   183 => (x"72",x"b2",x"73",x"4a"),
   184 => (x"26",x"4c",x"26",x"48"),
   185 => (x"26",x"4a",x"26",x"4b"),
   186 => (x"5a",x"5e",x"0e",x"4f"),
   187 => (x"0e",x"5d",x"5c",x"5b"),
   188 => (x"66",x"c4",x"8e",x"d0"),
   189 => (x"17",x"28",x"27",x"4c"),
   190 => (x"27",x"49",x"00",x"00"),
   191 => (x"00",x"00",x"17",x"30"),
   192 => (x"16",x"a8",x"27",x"79"),
   193 => (x"27",x"49",x"00",x"00"),
   194 => (x"00",x"00",x"16",x"f0"),
   195 => (x"16",x"f0",x"27",x"79"),
   196 => (x"27",x"49",x"00",x"00"),
   197 => (x"00",x"00",x"17",x"30"),
   198 => (x"16",x"f4",x"27",x"79"),
   199 => (x"c0",x"49",x"00",x"00"),
   200 => (x"16",x"f8",x"27",x"79"),
   201 => (x"c2",x"49",x"00",x"00"),
   202 => (x"16",x"fc",x"27",x"79"),
   203 => (x"c0",x"49",x"00",x"00"),
   204 => (x"00",x"27",x"79",x"e8"),
   205 => (x"49",x"00",x"00",x"17"),
   206 => (x"00",x"0f",x"fa",x"27"),
   207 => (x"1e",x"72",x"48",x"00"),
   208 => (x"10",x"4a",x"a1",x"df"),
   209 => (x"05",x"aa",x"71",x"51"),
   210 => (x"4a",x"26",x"87",x"f9"),
   211 => (x"00",x"16",x"b0",x"27"),
   212 => (x"19",x"27",x"49",x"00"),
   213 => (x"48",x"00",x"00",x"10"),
   214 => (x"a1",x"df",x"1e",x"72"),
   215 => (x"71",x"51",x"10",x"4a"),
   216 => (x"87",x"f9",x"05",x"aa"),
   217 => (x"9c",x"27",x"4a",x"26"),
   218 => (x"49",x"00",x"00",x"1e"),
   219 => (x"38",x"27",x"79",x"ca"),
   220 => (x"1e",x"00",x"00",x"10"),
   221 => (x"00",x"01",x"59",x"27"),
   222 => (x"86",x"c4",x"0f",x"00"),
   223 => (x"00",x"10",x"3a",x"27"),
   224 => (x"59",x"27",x"1e",x"00"),
   225 => (x"0f",x"00",x"00",x"01"),
   226 => (x"6a",x"27",x"86",x"c4"),
   227 => (x"1e",x"00",x"00",x"10"),
   228 => (x"00",x"01",x"59",x"27"),
   229 => (x"86",x"c4",x"0f",x"00"),
   230 => (x"00",x"16",x"1e",x"27"),
   231 => (x"c0",x"02",x"bf",x"00"),
   232 => (x"81",x"27",x"87",x"df"),
   233 => (x"1e",x"00",x"00",x"0e"),
   234 => (x"00",x"01",x"59",x"27"),
   235 => (x"86",x"c4",x"0f",x"00"),
   236 => (x"00",x"0e",x"ad",x"27"),
   237 => (x"59",x"27",x"1e",x"00"),
   238 => (x"0f",x"00",x"00",x"01"),
   239 => (x"dc",x"c0",x"86",x"c4"),
   240 => (x"0e",x"af",x"27",x"87"),
   241 => (x"27",x"1e",x"00",x"00"),
   242 => (x"00",x"00",x"01",x"59"),
   243 => (x"27",x"86",x"c4",x"0f"),
   244 => (x"00",x"00",x"0e",x"de"),
   245 => (x"01",x"59",x"27",x"1e"),
   246 => (x"c4",x"0f",x"00",x"00"),
   247 => (x"16",x"22",x"27",x"86"),
   248 => (x"1e",x"bf",x"00",x"00"),
   249 => (x"00",x"10",x"6c",x"27"),
   250 => (x"59",x"27",x"1e",x"00"),
   251 => (x"0f",x"00",x"00",x"01"),
   252 => (x"a5",x"27",x"86",x"c8"),
   253 => (x"0f",x"00",x"00",x"02"),
   254 => (x"a4",x"27",x"86",x"c0"),
   255 => (x"58",x"00",x"00",x"16"),
   256 => (x"22",x"27",x"4d",x"c1"),
   257 => (x"bf",x"00",x"00",x"16"),
   258 => (x"a9",x"b7",x"c0",x"49"),
   259 => (x"87",x"d7",x"c6",x"06"),
   260 => (x"00",x"0b",x"dc",x"27"),
   261 => (x"86",x"c0",x"0f",x"00"),
   262 => (x"00",x"0b",x"a0",x"27"),
   263 => (x"86",x"c0",x"0f",x"00"),
   264 => (x"79",x"c2",x"49",x"76"),
   265 => (x"d0",x"27",x"4c",x"c3"),
   266 => (x"49",x"00",x"00",x"16"),
   267 => (x"00",x"0e",x"ff",x"27"),
   268 => (x"1e",x"72",x"48",x"00"),
   269 => (x"10",x"4a",x"a1",x"df"),
   270 => (x"05",x"aa",x"71",x"51"),
   271 => (x"4a",x"26",x"87",x"f9"),
   272 => (x"c1",x"49",x"a6",x"c8"),
   273 => (x"16",x"d0",x"27",x"79"),
   274 => (x"1e",x"bf",x"00",x"00"),
   275 => (x"00",x"16",x"b0",x"27"),
   276 => (x"27",x"1e",x"bf",x"00"),
   277 => (x"00",x"00",x"0d",x"ab"),
   278 => (x"70",x"86",x"c8",x"0f"),
   279 => (x"05",x"9a",x"72",x"4a"),
   280 => (x"c1",x"87",x"c5",x"c0"),
   281 => (x"87",x"c2",x"c0",x"4a"),
   282 => (x"30",x"27",x"4a",x"c0"),
   283 => (x"49",x"00",x"00",x"18"),
   284 => (x"49",x"6e",x"79",x"72"),
   285 => (x"03",x"a9",x"b7",x"74"),
   286 => (x"6e",x"87",x"ed",x"c0"),
   287 => (x"72",x"92",x"c5",x"4a"),
   288 => (x"d0",x"88",x"74",x"48"),
   289 => (x"a6",x"cc",x"58",x"a6"),
   290 => (x"74",x"1e",x"72",x"4a"),
   291 => (x"1e",x"66",x"c8",x"1e"),
   292 => (x"00",x"0c",x"d0",x"27"),
   293 => (x"86",x"cc",x"0f",x"00"),
   294 => (x"80",x"c1",x"48",x"6e"),
   295 => (x"6e",x"58",x"a6",x"c4"),
   296 => (x"a9",x"b7",x"74",x"49"),
   297 => (x"87",x"d3",x"ff",x"04"),
   298 => (x"c4",x"1e",x"66",x"cc"),
   299 => (x"40",x"27",x"1e",x"66"),
   300 => (x"bf",x"00",x"00",x"18"),
   301 => (x"17",x"60",x"27",x"1e"),
   302 => (x"1e",x"bf",x"00",x"00"),
   303 => (x"00",x"0c",x"e5",x"27"),
   304 => (x"86",x"d0",x"0f",x"00"),
   305 => (x"00",x"16",x"a8",x"27"),
   306 => (x"27",x"1e",x"bf",x"00"),
   307 => (x"00",x"00",x"0a",x"8b"),
   308 => (x"c4",x"86",x"c4",x"0f"),
   309 => (x"c1",x"c1",x"49",x"a6"),
   310 => (x"18",x"28",x"27",x"51"),
   311 => (x"bf",x"97",x"00",x"00"),
   312 => (x"b7",x"32",x"d8",x"4a"),
   313 => (x"c1",x"49",x"72",x"2a"),
   314 => (x"04",x"a9",x"b7",x"c1"),
   315 => (x"c1",x"87",x"fb",x"c1"),
   316 => (x"c8",x"97",x"1e",x"c3"),
   317 => (x"32",x"d8",x"4a",x"66"),
   318 => (x"1e",x"72",x"2a",x"b7"),
   319 => (x"00",x"0d",x"73",x"27"),
   320 => (x"86",x"c8",x"0f",x"00"),
   321 => (x"66",x"c8",x"4a",x"70"),
   322 => (x"a9",x"b7",x"72",x"49"),
   323 => (x"87",x"f3",x"c0",x"05"),
   324 => (x"72",x"4a",x"a6",x"c8"),
   325 => (x"27",x"1e",x"c0",x"1e"),
   326 => (x"00",x"00",x"0c",x"51"),
   327 => (x"27",x"86",x"c8",x"0f"),
   328 => (x"00",x"00",x"16",x"d0"),
   329 => (x"0e",x"e0",x"27",x"49"),
   330 => (x"72",x"48",x"00",x"00"),
   331 => (x"4a",x"a1",x"df",x"1e"),
   332 => (x"aa",x"71",x"51",x"10"),
   333 => (x"26",x"87",x"f9",x"05"),
   334 => (x"27",x"4c",x"75",x"4a"),
   335 => (x"00",x"00",x"18",x"2c"),
   336 => (x"97",x"79",x"75",x"49"),
   337 => (x"c1",x"48",x"66",x"c4"),
   338 => (x"08",x"a6",x"c4",x"80"),
   339 => (x"66",x"c4",x"97",x"50"),
   340 => (x"b7",x"33",x"d8",x"4b"),
   341 => (x"18",x"28",x"27",x"2b"),
   342 => (x"bf",x"97",x"00",x"00"),
   343 => (x"b7",x"32",x"d8",x"4a"),
   344 => (x"72",x"49",x"73",x"2a"),
   345 => (x"fe",x"06",x"a9",x"b7"),
   346 => (x"94",x"6e",x"87",x"c5"),
   347 => (x"1e",x"72",x"49",x"74"),
   348 => (x"27",x"4a",x"66",x"d0"),
   349 => (x"00",x"00",x"0b",x"f0"),
   350 => (x"70",x"4a",x"26",x"0f"),
   351 => (x"58",x"a6",x"c4",x"48"),
   352 => (x"66",x"cc",x"4a",x"74"),
   353 => (x"72",x"92",x"c7",x"8a"),
   354 => (x"76",x"8c",x"6e",x"4c"),
   355 => (x"27",x"1e",x"72",x"4a"),
   356 => (x"00",x"00",x"0b",x"27"),
   357 => (x"c1",x"86",x"c4",x"0f"),
   358 => (x"27",x"49",x"75",x"85"),
   359 => (x"00",x"00",x"16",x"22"),
   360 => (x"06",x"a9",x"b7",x"bf"),
   361 => (x"27",x"87",x"e9",x"f9"),
   362 => (x"00",x"00",x"02",x"a5"),
   363 => (x"27",x"86",x"c0",x"0f"),
   364 => (x"00",x"00",x"17",x"24"),
   365 => (x"10",x"99",x"27",x"58"),
   366 => (x"27",x"1e",x"00",x"00"),
   367 => (x"00",x"00",x"01",x"59"),
   368 => (x"27",x"86",x"c4",x"0f"),
   369 => (x"00",x"00",x"10",x"a9"),
   370 => (x"01",x"59",x"27",x"1e"),
   371 => (x"c4",x"0f",x"00",x"00"),
   372 => (x"10",x"ab",x"27",x"86"),
   373 => (x"27",x"1e",x"00",x"00"),
   374 => (x"00",x"00",x"01",x"59"),
   375 => (x"27",x"86",x"c4",x"0f"),
   376 => (x"00",x"00",x"10",x"e1"),
   377 => (x"01",x"59",x"27",x"1e"),
   378 => (x"c4",x"0f",x"00",x"00"),
   379 => (x"18",x"2c",x"27",x"86"),
   380 => (x"1e",x"bf",x"00",x"00"),
   381 => (x"00",x"10",x"e3",x"27"),
   382 => (x"59",x"27",x"1e",x"00"),
   383 => (x"0f",x"00",x"00",x"01"),
   384 => (x"1e",x"c5",x"86",x"c8"),
   385 => (x"00",x"10",x"fc",x"27"),
   386 => (x"59",x"27",x"1e",x"00"),
   387 => (x"0f",x"00",x"00",x"01"),
   388 => (x"30",x"27",x"86",x"c8"),
   389 => (x"bf",x"00",x"00",x"18"),
   390 => (x"11",x"15",x"27",x"1e"),
   391 => (x"27",x"1e",x"00",x"00"),
   392 => (x"00",x"00",x"01",x"59"),
   393 => (x"c1",x"86",x"c8",x"0f"),
   394 => (x"11",x"2e",x"27",x"1e"),
   395 => (x"27",x"1e",x"00",x"00"),
   396 => (x"00",x"00",x"01",x"59"),
   397 => (x"27",x"86",x"c8",x"0f"),
   398 => (x"00",x"00",x"17",x"20"),
   399 => (x"d8",x"4a",x"bf",x"97"),
   400 => (x"72",x"2a",x"b7",x"32"),
   401 => (x"11",x"47",x"27",x"1e"),
   402 => (x"27",x"1e",x"00",x"00"),
   403 => (x"00",x"00",x"01",x"59"),
   404 => (x"c1",x"86",x"c8",x"0f"),
   405 => (x"60",x"27",x"1e",x"c1"),
   406 => (x"1e",x"00",x"00",x"11"),
   407 => (x"00",x"01",x"59",x"27"),
   408 => (x"86",x"c8",x"0f",x"00"),
   409 => (x"00",x"18",x"28",x"27"),
   410 => (x"4a",x"bf",x"97",x"00"),
   411 => (x"2a",x"b7",x"32",x"d8"),
   412 => (x"79",x"27",x"1e",x"72"),
   413 => (x"1e",x"00",x"00",x"11"),
   414 => (x"00",x"01",x"59",x"27"),
   415 => (x"86",x"c8",x"0f",x"00"),
   416 => (x"27",x"1e",x"c2",x"c1"),
   417 => (x"00",x"00",x"11",x"92"),
   418 => (x"01",x"59",x"27",x"1e"),
   419 => (x"c8",x"0f",x"00",x"00"),
   420 => (x"17",x"80",x"27",x"86"),
   421 => (x"1e",x"bf",x"00",x"00"),
   422 => (x"00",x"11",x"ab",x"27"),
   423 => (x"59",x"27",x"1e",x"00"),
   424 => (x"0f",x"00",x"00",x"01"),
   425 => (x"1e",x"c7",x"86",x"c8"),
   426 => (x"00",x"11",x"c4",x"27"),
   427 => (x"59",x"27",x"1e",x"00"),
   428 => (x"0f",x"00",x"00",x"01"),
   429 => (x"9c",x"27",x"86",x"c8"),
   430 => (x"bf",x"00",x"00",x"1e"),
   431 => (x"11",x"dd",x"27",x"1e"),
   432 => (x"27",x"1e",x"00",x"00"),
   433 => (x"00",x"00",x"01",x"59"),
   434 => (x"27",x"86",x"c8",x"0f"),
   435 => (x"00",x"00",x"11",x"f6"),
   436 => (x"01",x"59",x"27",x"1e"),
   437 => (x"c4",x"0f",x"00",x"00"),
   438 => (x"12",x"20",x"27",x"86"),
   439 => (x"27",x"1e",x"00",x"00"),
   440 => (x"00",x"00",x"01",x"59"),
   441 => (x"a8",x"86",x"c4",x"0f"),
   442 => (x"bf",x"00",x"00",x"16"),
   443 => (x"12",x"2c",x"27",x"1e"),
   444 => (x"27",x"1e",x"00",x"00"),
   445 => (x"00",x"00",x"01",x"59"),
   446 => (x"27",x"86",x"c8",x"0f"),
   447 => (x"00",x"00",x"12",x"45"),
   448 => (x"01",x"59",x"27",x"1e"),
   449 => (x"c4",x"0f",x"00",x"00"),
   450 => (x"16",x"a8",x"27",x"86"),
   451 => (x"4a",x"bf",x"00",x"00"),
   452 => (x"1e",x"6a",x"82",x"c4"),
   453 => (x"00",x"12",x"76",x"27"),
   454 => (x"59",x"27",x"1e",x"00"),
   455 => (x"0f",x"00",x"00",x"01"),
   456 => (x"1e",x"c0",x"86",x"c8"),
   457 => (x"00",x"12",x"8f",x"27"),
   458 => (x"59",x"27",x"1e",x"00"),
   459 => (x"0f",x"00",x"00",x"01"),
   460 => (x"a8",x"27",x"86",x"c8"),
   461 => (x"bf",x"00",x"00",x"16"),
   462 => (x"6a",x"82",x"c8",x"4a"),
   463 => (x"12",x"a8",x"27",x"1e"),
   464 => (x"27",x"1e",x"00",x"00"),
   465 => (x"00",x"00",x"01",x"59"),
   466 => (x"c2",x"86",x"c8",x"0f"),
   467 => (x"12",x"c1",x"27",x"1e"),
   468 => (x"27",x"1e",x"00",x"00"),
   469 => (x"00",x"00",x"01",x"59"),
   470 => (x"27",x"86",x"c8",x"0f"),
   471 => (x"00",x"00",x"16",x"a8"),
   472 => (x"82",x"cc",x"4a",x"bf"),
   473 => (x"da",x"27",x"1e",x"6a"),
   474 => (x"1e",x"00",x"00",x"12"),
   475 => (x"00",x"01",x"59",x"27"),
   476 => (x"86",x"c8",x"0f",x"00"),
   477 => (x"f3",x"27",x"1e",x"d1"),
   478 => (x"1e",x"00",x"00",x"12"),
   479 => (x"00",x"01",x"59",x"27"),
   480 => (x"86",x"c8",x"0f",x"00"),
   481 => (x"00",x"16",x"a8",x"27"),
   482 => (x"d0",x"4a",x"bf",x"00"),
   483 => (x"27",x"1e",x"72",x"82"),
   484 => (x"00",x"00",x"13",x"0c"),
   485 => (x"01",x"59",x"27",x"1e"),
   486 => (x"c8",x"0f",x"00",x"00"),
   487 => (x"13",x"25",x"27",x"86"),
   488 => (x"27",x"1e",x"00",x"00"),
   489 => (x"00",x"00",x"01",x"59"),
   490 => (x"27",x"86",x"c4",x"0f"),
   491 => (x"00",x"00",x"13",x"5a"),
   492 => (x"01",x"59",x"27",x"1e"),
   493 => (x"c4",x"0f",x"00",x"00"),
   494 => (x"00",x"17",x"28",x"86"),
   495 => (x"27",x"1e",x"bf",x"00"),
   496 => (x"00",x"00",x"13",x"6b"),
   497 => (x"01",x"59",x"27",x"1e"),
   498 => (x"c8",x"0f",x"00",x"00"),
   499 => (x"13",x"84",x"27",x"86"),
   500 => (x"27",x"1e",x"00",x"00"),
   501 => (x"00",x"00",x"01",x"59"),
   502 => (x"27",x"86",x"c4",x"0f"),
   503 => (x"00",x"00",x"17",x"28"),
   504 => (x"82",x"c4",x"4a",x"bf"),
   505 => (x"c4",x"27",x"1e",x"6a"),
   506 => (x"1e",x"00",x"00",x"13"),
   507 => (x"00",x"01",x"59",x"27"),
   508 => (x"86",x"c8",x"0f",x"00"),
   509 => (x"dd",x"27",x"1e",x"c0"),
   510 => (x"1e",x"00",x"00",x"13"),
   511 => (x"00",x"01",x"59",x"27"),
   512 => (x"86",x"c8",x"0f",x"00"),
   513 => (x"00",x"17",x"28",x"27"),
   514 => (x"c8",x"4a",x"bf",x"00"),
   515 => (x"27",x"1e",x"6a",x"82"),
   516 => (x"00",x"00",x"13",x"f6"),
   517 => (x"01",x"59",x"27",x"1e"),
   518 => (x"c8",x"0f",x"00",x"00"),
   519 => (x"27",x"1e",x"c1",x"86"),
   520 => (x"00",x"00",x"14",x"0f"),
   521 => (x"01",x"59",x"27",x"1e"),
   522 => (x"c8",x"0f",x"00",x"00"),
   523 => (x"17",x"28",x"27",x"86"),
   524 => (x"4a",x"bf",x"00",x"00"),
   525 => (x"1e",x"6a",x"82",x"cc"),
   526 => (x"00",x"14",x"28",x"27"),
   527 => (x"59",x"27",x"1e",x"00"),
   528 => (x"0f",x"00",x"00",x"01"),
   529 => (x"1e",x"d2",x"86",x"c8"),
   530 => (x"00",x"14",x"41",x"27"),
   531 => (x"59",x"27",x"1e",x"00"),
   532 => (x"0f",x"00",x"00",x"01"),
   533 => (x"28",x"27",x"86",x"c8"),
   534 => (x"bf",x"00",x"00",x"17"),
   535 => (x"72",x"82",x"d0",x"4a"),
   536 => (x"14",x"5a",x"27",x"1e"),
   537 => (x"27",x"1e",x"00",x"00"),
   538 => (x"00",x"00",x"01",x"59"),
   539 => (x"27",x"86",x"c8",x"0f"),
   540 => (x"00",x"00",x"14",x"73"),
   541 => (x"01",x"59",x"27",x"1e"),
   542 => (x"c4",x"0f",x"00",x"00"),
   543 => (x"27",x"1e",x"6e",x"86"),
   544 => (x"00",x"00",x"14",x"a8"),
   545 => (x"01",x"59",x"27",x"1e"),
   546 => (x"c8",x"0f",x"00",x"00"),
   547 => (x"27",x"1e",x"c5",x"86"),
   548 => (x"00",x"00",x"14",x"c1"),
   549 => (x"01",x"59",x"27",x"1e"),
   550 => (x"c8",x"0f",x"00",x"00"),
   551 => (x"27",x"1e",x"74",x"86"),
   552 => (x"00",x"00",x"14",x"da"),
   553 => (x"01",x"59",x"27",x"1e"),
   554 => (x"c8",x"0f",x"00",x"00"),
   555 => (x"27",x"1e",x"cd",x"86"),
   556 => (x"00",x"00",x"14",x"f3"),
   557 => (x"01",x"59",x"27",x"1e"),
   558 => (x"c8",x"0f",x"00",x"00"),
   559 => (x"1e",x"66",x"cc",x"86"),
   560 => (x"00",x"15",x"0c",x"27"),
   561 => (x"59",x"27",x"1e",x"00"),
   562 => (x"0f",x"00",x"00",x"01"),
   563 => (x"1e",x"c7",x"86",x"c8"),
   564 => (x"00",x"15",x"25",x"27"),
   565 => (x"59",x"27",x"1e",x"00"),
   566 => (x"0f",x"00",x"00",x"01"),
   567 => (x"66",x"c8",x"86",x"c8"),
   568 => (x"15",x"3e",x"27",x"1e"),
   569 => (x"27",x"1e",x"00",x"00"),
   570 => (x"00",x"00",x"01",x"59"),
   571 => (x"c1",x"86",x"c8",x"0f"),
   572 => (x"15",x"57",x"27",x"1e"),
   573 => (x"27",x"1e",x"00",x"00"),
   574 => (x"00",x"00",x"01",x"59"),
   575 => (x"27",x"86",x"c8",x"0f"),
   576 => (x"00",x"00",x"16",x"b0"),
   577 => (x"70",x"27",x"1e",x"bf"),
   578 => (x"1e",x"00",x"00",x"15"),
   579 => (x"00",x"01",x"59",x"27"),
   580 => (x"86",x"c8",x"0f",x"00"),
   581 => (x"00",x"15",x"89",x"27"),
   582 => (x"59",x"27",x"1e",x"00"),
   583 => (x"0f",x"00",x"00",x"01"),
   584 => (x"d0",x"27",x"86",x"c4"),
   585 => (x"bf",x"00",x"00",x"16"),
   586 => (x"15",x"be",x"27",x"1e"),
   587 => (x"27",x"1e",x"00",x"00"),
   588 => (x"00",x"00",x"01",x"59"),
   589 => (x"27",x"86",x"c8",x"0f"),
   590 => (x"00",x"00",x"15",x"d7"),
   591 => (x"01",x"59",x"27",x"1e"),
   592 => (x"c4",x"0f",x"00",x"00"),
   593 => (x"16",x"0c",x"27",x"86"),
   594 => (x"27",x"1e",x"00",x"00"),
   595 => (x"00",x"00",x"01",x"59"),
   596 => (x"27",x"86",x"c4",x"0f"),
   597 => (x"00",x"00",x"17",x"24"),
   598 => (x"a4",x"27",x"4a",x"bf"),
   599 => (x"bf",x"00",x"00",x"16"),
   600 => (x"16",x"ac",x"27",x"8a"),
   601 => (x"72",x"49",x"00",x"00"),
   602 => (x"27",x"1e",x"72",x"79"),
   603 => (x"00",x"00",x"16",x"0e"),
   604 => (x"01",x"59",x"27",x"1e"),
   605 => (x"c8",x"0f",x"00",x"00"),
   606 => (x"16",x"ac",x"27",x"86"),
   607 => (x"49",x"bf",x"00",x"00"),
   608 => (x"a9",x"b7",x"f8",x"c1"),
   609 => (x"87",x"ea",x"c0",x"03"),
   610 => (x"00",x"0f",x"1e",x"27"),
   611 => (x"59",x"27",x"1e",x"00"),
   612 => (x"0f",x"00",x"00",x"01"),
   613 => (x"54",x"27",x"86",x"c4"),
   614 => (x"1e",x"00",x"00",x"0f"),
   615 => (x"00",x"01",x"59",x"27"),
   616 => (x"86",x"c4",x"0f",x"00"),
   617 => (x"00",x"0f",x"74",x"27"),
   618 => (x"59",x"27",x"1e",x"00"),
   619 => (x"0f",x"00",x"00",x"01"),
   620 => (x"ac",x"27",x"86",x"c4"),
   621 => (x"bf",x"00",x"00",x"16"),
   622 => (x"cf",x"4b",x"72",x"4a"),
   623 => (x"49",x"73",x"93",x"e8"),
   624 => (x"22",x"27",x"1e",x"72"),
   625 => (x"bf",x"00",x"00",x"16"),
   626 => (x"0b",x"f0",x"27",x"4a"),
   627 => (x"26",x"0f",x"00",x"00"),
   628 => (x"27",x"48",x"70",x"4a"),
   629 => (x"00",x"00",x"17",x"2c"),
   630 => (x"16",x"22",x"27",x"58"),
   631 => (x"4b",x"bf",x"00",x"00"),
   632 => (x"e8",x"cf",x"4c",x"73"),
   633 => (x"72",x"49",x"74",x"94"),
   634 => (x"27",x"4a",x"72",x"1e"),
   635 => (x"00",x"00",x"0b",x"f0"),
   636 => (x"70",x"4a",x"26",x"0f"),
   637 => (x"16",x"a0",x"27",x"48"),
   638 => (x"c8",x"58",x"00",x"00"),
   639 => (x"49",x"73",x"93",x"f9"),
   640 => (x"4a",x"72",x"1e",x"72"),
   641 => (x"00",x"0b",x"f0",x"27"),
   642 => (x"4a",x"26",x"0f",x"00"),
   643 => (x"34",x"27",x"48",x"70"),
   644 => (x"58",x"00",x"00",x"18"),
   645 => (x"00",x"0f",x"76",x"27"),
   646 => (x"59",x"27",x"1e",x"00"),
   647 => (x"0f",x"00",x"00",x"01"),
   648 => (x"2c",x"27",x"86",x"c4"),
   649 => (x"bf",x"00",x"00",x"17"),
   650 => (x"0f",x"a3",x"27",x"1e"),
   651 => (x"27",x"1e",x"00",x"00"),
   652 => (x"00",x"00",x"01",x"59"),
   653 => (x"27",x"86",x"c8",x"0f"),
   654 => (x"00",x"00",x"0f",x"a8"),
   655 => (x"01",x"59",x"27",x"1e"),
   656 => (x"c4",x"0f",x"00",x"00"),
   657 => (x"16",x"a0",x"27",x"86"),
   658 => (x"1e",x"bf",x"00",x"00"),
   659 => (x"00",x"0f",x"d5",x"27"),
   660 => (x"59",x"27",x"1e",x"00"),
   661 => (x"0f",x"00",x"00",x"01"),
   662 => (x"34",x"27",x"86",x"c8"),
   663 => (x"bf",x"00",x"00",x"18"),
   664 => (x"0f",x"da",x"27",x"1e"),
   665 => (x"27",x"1e",x"00",x"00"),
   666 => (x"00",x"00",x"01",x"59"),
   667 => (x"27",x"86",x"c8",x"0f"),
   668 => (x"00",x"00",x"0f",x"f8"),
   669 => (x"01",x"59",x"27",x"1e"),
   670 => (x"c4",x"0f",x"00",x"00"),
   671 => (x"d0",x"48",x"c0",x"86"),
   672 => (x"26",x"4d",x"26",x"86"),
   673 => (x"26",x"4b",x"26",x"4c"),
   674 => (x"0e",x"4f",x"26",x"4a"),
   675 => (x"5c",x"5b",x"5a",x"5e"),
   676 => (x"a6",x"d4",x"0e",x"5d"),
   677 => (x"72",x"4a",x"bf",x"bf"),
   678 => (x"00",x"16",x"a8",x"4d"),
   679 => (x"72",x"48",x"bf",x"00"),
   680 => (x"a1",x"f0",x"c0",x"1e"),
   681 => (x"71",x"51",x"10",x"4a"),
   682 => (x"87",x"f9",x"05",x"aa"),
   683 => (x"66",x"d4",x"4a",x"26"),
   684 => (x"c5",x"84",x"cc",x"4c"),
   685 => (x"cc",x"4b",x"72",x"7c"),
   686 => (x"d4",x"7b",x"6c",x"83"),
   687 => (x"7a",x"bf",x"bf",x"a6"),
   688 => (x"69",x"27",x"1e",x"72"),
   689 => (x"0f",x"00",x"00",x"0b"),
   690 => (x"82",x"c4",x"86",x"c4"),
   691 => (x"c0",x"05",x"9a",x"6a"),
   692 => (x"4b",x"75",x"87",x"f2"),
   693 => (x"4a",x"75",x"83",x"c8"),
   694 => (x"7a",x"c6",x"82",x"cc"),
   695 => (x"66",x"d8",x"1e",x"73"),
   696 => (x"6b",x"83",x"c8",x"4b"),
   697 => (x"0c",x"51",x"27",x"1e"),
   698 => (x"c8",x"0f",x"00",x"00"),
   699 => (x"00",x"16",x"a8",x"86"),
   700 => (x"72",x"7d",x"bf",x"00"),
   701 => (x"6a",x"1e",x"ca",x"1e"),
   702 => (x"0c",x"d0",x"27",x"1e"),
   703 => (x"cc",x"0f",x"00",x"00"),
   704 => (x"87",x"d9",x"c0",x"86"),
   705 => (x"bf",x"bf",x"a6",x"d4"),
   706 => (x"bf",x"a6",x"d4",x"4a"),
   707 => (x"1e",x"72",x"48",x"49"),
   708 => (x"4a",x"a1",x"f0",x"c0"),
   709 => (x"aa",x"71",x"51",x"10"),
   710 => (x"26",x"87",x"f9",x"05"),
   711 => (x"26",x"4d",x"26",x"4a"),
   712 => (x"26",x"4b",x"26",x"4c"),
   713 => (x"0e",x"4f",x"26",x"4a"),
   714 => (x"0e",x"5b",x"5a",x"5e"),
   715 => (x"bf",x"a6",x"d0",x"1e"),
   716 => (x"83",x"ca",x"4b",x"bf"),
   717 => (x"00",x"17",x"20",x"27"),
   718 => (x"4a",x"bf",x"97",x"00"),
   719 => (x"2a",x"b7",x"32",x"d8"),
   720 => (x"c1",x"c1",x"49",x"72"),
   721 => (x"c0",x"05",x"a9",x"b7"),
   722 => (x"8b",x"c1",x"87",x"d3"),
   723 => (x"2c",x"27",x"48",x"73"),
   724 => (x"bf",x"00",x"00",x"18"),
   725 => (x"49",x"66",x"d0",x"88"),
   726 => (x"c0",x"49",x"76",x"58"),
   727 => (x"ff",x"05",x"6e",x"79"),
   728 => (x"26",x"26",x"87",x"d2"),
   729 => (x"26",x"4a",x"26",x"4b"),
   730 => (x"1e",x"72",x"1e",x"4f"),
   731 => (x"00",x"16",x"a8",x"27"),
   732 => (x"c0",x"02",x"bf",x"00"),
   733 => (x"a6",x"c8",x"87",x"ca"),
   734 => (x"16",x"a8",x"49",x"bf"),
   735 => (x"79",x"bf",x"00",x"00"),
   736 => (x"00",x"16",x"a8",x"27"),
   737 => (x"cc",x"4a",x"bf",x"00"),
   738 => (x"27",x"1e",x"72",x"82"),
   739 => (x"00",x"00",x"18",x"2c"),
   740 => (x"1e",x"ca",x"1e",x"bf"),
   741 => (x"00",x"0c",x"d0",x"27"),
   742 => (x"86",x"cc",x"0f",x"00"),
   743 => (x"4f",x"26",x"4a",x"26"),
   744 => (x"27",x"1e",x"72",x"1e"),
   745 => (x"00",x"00",x"17",x"20"),
   746 => (x"d8",x"4a",x"bf",x"97"),
   747 => (x"72",x"2a",x"b7",x"32"),
   748 => (x"b7",x"c1",x"c1",x"49"),
   749 => (x"c5",x"c0",x"02",x"a9"),
   750 => (x"c0",x"4a",x"c0",x"87"),
   751 => (x"4a",x"c1",x"87",x"c2"),
   752 => (x"00",x"18",x"30",x"27"),
   753 => (x"72",x"48",x"bf",x"00"),
   754 => (x"18",x"30",x"27",x"b0"),
   755 => (x"27",x"58",x"00",x"00"),
   756 => (x"00",x"00",x"18",x"28"),
   757 => (x"51",x"c2",x"c1",x"49"),
   758 => (x"4f",x"26",x"4a",x"26"),
   759 => (x"17",x"20",x"27",x"1e"),
   760 => (x"c1",x"49",x"00",x"00"),
   761 => (x"30",x"27",x"51",x"c1"),
   762 => (x"49",x"00",x"00",x"18"),
   763 => (x"4f",x"26",x"79",x"c0"),
   764 => (x"72",x"1e",x"73",x"1e"),
   765 => (x"87",x"d9",x"02",x"9a"),
   766 => (x"4b",x"c1",x"48",x"c0"),
   767 => (x"82",x"01",x"a9",x"72"),
   768 => (x"87",x"f8",x"83",x"73"),
   769 => (x"89",x"03",x"a9",x"72"),
   770 => (x"c1",x"07",x"80",x"73"),
   771 => (x"f3",x"05",x"2b",x"2a"),
   772 => (x"26",x"4b",x"26",x"87"),
   773 => (x"1e",x"75",x"1e",x"4f"),
   774 => (x"a1",x"71",x"4d",x"c0"),
   775 => (x"c1",x"b9",x"ff",x"04"),
   776 => (x"72",x"07",x"bd",x"81"),
   777 => (x"ba",x"ff",x"04",x"a2"),
   778 => (x"07",x"bd",x"82",x"c1"),
   779 => (x"9d",x"75",x"87",x"c2"),
   780 => (x"c1",x"b8",x"ff",x"05"),
   781 => (x"4d",x"25",x"07",x"80"),
   782 => (x"72",x"1e",x"4f",x"26"),
   783 => (x"49",x"66",x"c8",x"1e"),
   784 => (x"11",x"4a",x"66",x"cc"),
   785 => (x"c4",x"02",x"12",x"48"),
   786 => (x"f6",x"02",x"88",x"87"),
   787 => (x"26",x"4a",x"26",x"87"),
   788 => (x"5a",x"5e",x"0e",x"4f"),
   789 => (x"66",x"d0",x"0e",x"5b"),
   790 => (x"7b",x"66",x"cc",x"4b"),
   791 => (x"27",x"1e",x"66",x"cc"),
   792 => (x"00",x"00",x"0e",x"5c"),
   793 => (x"70",x"86",x"c4",x"0f"),
   794 => (x"05",x"9a",x"72",x"4a"),
   795 => (x"c3",x"87",x"c2",x"c0"),
   796 => (x"4a",x"66",x"cc",x"7b"),
   797 => (x"c0",x"49",x"66",x"cc"),
   798 => (x"c0",x"02",x"a9",x"b7"),
   799 => (x"49",x"72",x"87",x"e7"),
   800 => (x"02",x"a9",x"b7",x"c1"),
   801 => (x"72",x"87",x"e3",x"c0"),
   802 => (x"a9",x"b7",x"c2",x"49"),
   803 => (x"87",x"f3",x"c0",x"02"),
   804 => (x"b7",x"c3",x"49",x"72"),
   805 => (x"f1",x"c0",x"02",x"a9"),
   806 => (x"c4",x"49",x"72",x"87"),
   807 => (x"c0",x"02",x"a9",x"b7"),
   808 => (x"e5",x"c0",x"87",x"e6"),
   809 => (x"c0",x"7b",x"c0",x"87"),
   810 => (x"2c",x"27",x"87",x"e0"),
   811 => (x"bf",x"00",x"00",x"18"),
   812 => (x"b7",x"e4",x"c1",x"49"),
   813 => (x"c5",x"c0",x"06",x"a9"),
   814 => (x"c0",x"7b",x"c0",x"87"),
   815 => (x"7b",x"c3",x"87",x"cc"),
   816 => (x"c1",x"87",x"c7",x"c0"),
   817 => (x"87",x"c2",x"c0",x"7b"),
   818 => (x"4b",x"26",x"7b",x"c2"),
   819 => (x"4f",x"26",x"4a",x"26"),
   820 => (x"c8",x"1e",x"72",x"1e"),
   821 => (x"82",x"c2",x"4a",x"66"),
   822 => (x"72",x"48",x"66",x"cc"),
   823 => (x"49",x"66",x"d0",x"80"),
   824 => (x"26",x"4a",x"26",x"58"),
   825 => (x"5a",x"5e",x"0e",x"4f"),
   826 => (x"0e",x"5d",x"5c",x"5b"),
   827 => (x"c5",x"4d",x"66",x"dc"),
   828 => (x"c4",x"4a",x"75",x"85"),
   829 => (x"d4",x"4a",x"72",x"92"),
   830 => (x"e0",x"c0",x"82",x"66"),
   831 => (x"4b",x"72",x"7a",x"66"),
   832 => (x"7b",x"6a",x"83",x"c4"),
   833 => (x"75",x"82",x"f8",x"c1"),
   834 => (x"75",x"4c",x"75",x"7a"),
   835 => (x"75",x"82",x"c1",x"4a"),
   836 => (x"a9",x"b7",x"72",x"49"),
   837 => (x"87",x"e3",x"c0",x"01"),
   838 => (x"c8",x"c3",x"4b",x"75"),
   839 => (x"d8",x"4b",x"73",x"93"),
   840 => (x"4a",x"74",x"83",x"66"),
   841 => (x"4a",x"72",x"92",x"c4"),
   842 => (x"7a",x"75",x"82",x"73"),
   843 => (x"4a",x"75",x"84",x"c1"),
   844 => (x"49",x"74",x"82",x"c1"),
   845 => (x"06",x"a9",x"b7",x"72"),
   846 => (x"75",x"87",x"dd",x"ff"),
   847 => (x"94",x"c8",x"c3",x"4c"),
   848 => (x"66",x"d8",x"4c",x"74"),
   849 => (x"c4",x"4a",x"75",x"84"),
   850 => (x"72",x"4b",x"74",x"92"),
   851 => (x"c1",x"48",x"6b",x"83"),
   852 => (x"66",x"d4",x"58",x"80"),
   853 => (x"c0",x"83",x"72",x"4b"),
   854 => (x"72",x"84",x"e0",x"fe"),
   855 => (x"6b",x"82",x"74",x"4a"),
   856 => (x"18",x"2c",x"27",x"7a"),
   857 => (x"c5",x"49",x"00",x"00"),
   858 => (x"26",x"4d",x"26",x"79"),
   859 => (x"26",x"4b",x"26",x"4c"),
   860 => (x"0e",x"4f",x"26",x"4a"),
   861 => (x"5c",x"5b",x"5a",x"5e"),
   862 => (x"66",x"d0",x"97",x"0e"),
   863 => (x"d8",x"4b",x"74",x"4c"),
   864 => (x"97",x"2b",x"b7",x"33"),
   865 => (x"d8",x"4a",x"66",x"d4"),
   866 => (x"73",x"2a",x"b7",x"32"),
   867 => (x"a9",x"b7",x"72",x"49"),
   868 => (x"87",x"c5",x"c0",x"02"),
   869 => (x"ca",x"c0",x"48",x"c0"),
   870 => (x"17",x"20",x"27",x"87"),
   871 => (x"74",x"49",x"00",x"00"),
   872 => (x"26",x"48",x"c1",x"51"),
   873 => (x"26",x"4b",x"26",x"4c"),
   874 => (x"0e",x"4f",x"26",x"4a"),
   875 => (x"0e",x"5b",x"5a",x"5e"),
   876 => (x"d4",x"4b",x"c2",x"1e"),
   877 => (x"82",x"c1",x"4a",x"66"),
   878 => (x"6a",x"97",x"82",x"73"),
   879 => (x"b7",x"32",x"d8",x"4a"),
   880 => (x"d4",x"1e",x"72",x"2a"),
   881 => (x"82",x"73",x"4a",x"66"),
   882 => (x"d8",x"4a",x"6a",x"97"),
   883 => (x"72",x"2a",x"b7",x"32"),
   884 => (x"0d",x"73",x"27",x"1e"),
   885 => (x"c8",x"0f",x"00",x"00"),
   886 => (x"72",x"4a",x"70",x"86"),
   887 => (x"c7",x"c0",x"05",x"9a"),
   888 => (x"c1",x"49",x"76",x"87"),
   889 => (x"83",x"c1",x"51",x"c1"),
   890 => (x"b7",x"c2",x"49",x"73"),
   891 => (x"c2",x"ff",x"06",x"a9"),
   892 => (x"4a",x"6e",x"97",x"87"),
   893 => (x"2a",x"b7",x"32",x"d8"),
   894 => (x"d7",x"c1",x"49",x"72"),
   895 => (x"c0",x"04",x"a9",x"b7"),
   896 => (x"6e",x"97",x"87",x"d3"),
   897 => (x"b7",x"32",x"d8",x"4a"),
   898 => (x"c1",x"49",x"72",x"2a"),
   899 => (x"03",x"a9",x"b7",x"da"),
   900 => (x"c7",x"87",x"c2",x"c0"),
   901 => (x"4a",x"6e",x"97",x"4b"),
   902 => (x"2a",x"b7",x"32",x"d8"),
   903 => (x"d2",x"c1",x"49",x"72"),
   904 => (x"c0",x"05",x"a9",x"b7"),
   905 => (x"48",x"c1",x"87",x"c5"),
   906 => (x"d4",x"87",x"ea",x"c0"),
   907 => (x"66",x"d4",x"1e",x"66"),
   908 => (x"0c",x"3a",x"27",x"1e"),
   909 => (x"c8",x"0f",x"00",x"00"),
   910 => (x"72",x"4a",x"70",x"86"),
   911 => (x"a9",x"b7",x"c0",x"49"),
   912 => (x"87",x"cf",x"c0",x"06"),
   913 => (x"80",x"c7",x"48",x"73"),
   914 => (x"00",x"18",x"2c",x"27"),
   915 => (x"48",x"c1",x"58",x"00"),
   916 => (x"c0",x"87",x"c2",x"c0"),
   917 => (x"4b",x"26",x"26",x"48"),
   918 => (x"4f",x"26",x"4a",x"26"),
   919 => (x"49",x"66",x"c4",x"1e"),
   920 => (x"05",x"a9",x"b7",x"c2"),
   921 => (x"c1",x"87",x"c5",x"c0"),
   922 => (x"87",x"c2",x"c0",x"48"),
   923 => (x"4f",x"26",x"48",x"c0"),
   924 => (x"33",x"32",x"31",x"30"),
   925 => (x"37",x"36",x"35",x"34"),
   926 => (x"42",x"41",x"39",x"38"),
   927 => (x"46",x"45",x"44",x"43"),
   928 => (x"6f",x"72",x"50",x"00"),
   929 => (x"6d",x"61",x"72",x"67"),
   930 => (x"6d",x"6f",x"63",x"20"),
   931 => (x"65",x"6c",x"69",x"70"),
   932 => (x"69",x"77",x"20",x"64"),
   933 => (x"27",x"20",x"68",x"74"),
   934 => (x"69",x"67",x"65",x"72"),
   935 => (x"72",x"65",x"74",x"73"),
   936 => (x"74",x"61",x"20",x"27"),
   937 => (x"62",x"69",x"72",x"74"),
   938 => (x"0a",x"65",x"74",x"75"),
   939 => (x"50",x"00",x"0a",x"00"),
   940 => (x"72",x"67",x"6f",x"72"),
   941 => (x"63",x"20",x"6d",x"61"),
   942 => (x"69",x"70",x"6d",x"6f"),
   943 => (x"20",x"64",x"65",x"6c"),
   944 => (x"68",x"74",x"69",x"77"),
   945 => (x"20",x"74",x"75",x"6f"),
   946 => (x"67",x"65",x"72",x"27"),
   947 => (x"65",x"74",x"73",x"69"),
   948 => (x"61",x"20",x"27",x"72"),
   949 => (x"69",x"72",x"74",x"74"),
   950 => (x"65",x"74",x"75",x"62"),
   951 => (x"00",x"0a",x"00",x"0a"),
   952 => (x"59",x"52",x"48",x"44"),
   953 => (x"4e",x"4f",x"54",x"53"),
   954 => (x"52",x"50",x"20",x"45"),
   955 => (x"41",x"52",x"47",x"4f"),
   956 => (x"33",x"20",x"2c",x"4d"),
   957 => (x"20",x"44",x"52",x"27"),
   958 => (x"49",x"52",x"54",x"53"),
   959 => (x"44",x"00",x"47",x"4e"),
   960 => (x"53",x"59",x"52",x"48"),
   961 => (x"45",x"4e",x"4f",x"54"),
   962 => (x"4f",x"52",x"50",x"20"),
   963 => (x"4d",x"41",x"52",x"47"),
   964 => (x"27",x"32",x"20",x"2c"),
   965 => (x"53",x"20",x"44",x"4e"),
   966 => (x"4e",x"49",x"52",x"54"),
   967 => (x"65",x"4d",x"00",x"47"),
   968 => (x"72",x"75",x"73",x"61"),
   969 => (x"74",x"20",x"64",x"65"),
   970 => (x"20",x"65",x"6d",x"69"),
   971 => (x"20",x"6f",x"6f",x"74"),
   972 => (x"6c",x"61",x"6d",x"73"),
   973 => (x"6f",x"74",x"20",x"6c"),
   974 => (x"74",x"62",x"6f",x"20"),
   975 => (x"20",x"6e",x"69",x"61"),
   976 => (x"6e",x"61",x"65",x"6d"),
   977 => (x"66",x"67",x"6e",x"69"),
   978 => (x"72",x"20",x"6c",x"75"),
   979 => (x"6c",x"75",x"73",x"65"),
   980 => (x"00",x"0a",x"73",x"74"),
   981 => (x"61",x"65",x"6c",x"50"),
   982 => (x"69",x"20",x"65",x"73"),
   983 => (x"65",x"72",x"63",x"6e"),
   984 => (x"20",x"65",x"73",x"61"),
   985 => (x"62",x"6d",x"75",x"6e"),
   986 => (x"6f",x"20",x"72",x"65"),
   987 => (x"75",x"72",x"20",x"66"),
   988 => (x"00",x"0a",x"73",x"6e"),
   989 => (x"69",x"4d",x"00",x"0a"),
   990 => (x"73",x"6f",x"72",x"63"),
   991 => (x"6e",x"6f",x"63",x"65"),
   992 => (x"66",x"20",x"73",x"64"),
   993 => (x"6f",x"20",x"72",x"6f"),
   994 => (x"72",x"20",x"65",x"6e"),
   995 => (x"74",x"20",x"6e",x"75"),
   996 => (x"75",x"6f",x"72",x"68"),
   997 => (x"44",x"20",x"68",x"67"),
   998 => (x"73",x"79",x"72",x"68"),
   999 => (x"65",x"6e",x"6f",x"74"),
  1000 => (x"25",x"00",x"20",x"3a"),
  1001 => (x"00",x"0a",x"20",x"64"),
  1002 => (x"79",x"72",x"68",x"44"),
  1003 => (x"6e",x"6f",x"74",x"73"),
  1004 => (x"70",x"20",x"73",x"65"),
  1005 => (x"53",x"20",x"72",x"65"),
  1006 => (x"6e",x"6f",x"63",x"65"),
  1007 => (x"20",x"20",x"3a",x"64"),
  1008 => (x"20",x"20",x"20",x"20"),
  1009 => (x"20",x"20",x"20",x"20"),
  1010 => (x"20",x"20",x"20",x"20"),
  1011 => (x"20",x"20",x"20",x"20"),
  1012 => (x"20",x"20",x"20",x"20"),
  1013 => (x"20",x"64",x"25",x"00"),
  1014 => (x"41",x"56",x"00",x"0a"),
  1015 => (x"49",x"4d",x"20",x"58"),
  1016 => (x"72",x"20",x"53",x"50"),
  1017 => (x"6e",x"69",x"74",x"61"),
  1018 => (x"20",x"2a",x"20",x"67"),
  1019 => (x"30",x"30",x"30",x"31"),
  1020 => (x"25",x"20",x"3d",x"20"),
  1021 => (x"00",x"0a",x"20",x"64"),
  1022 => (x"48",x"44",x"00",x"0a"),
  1023 => (x"54",x"53",x"59",x"52"),
  1024 => (x"20",x"45",x"4e",x"4f"),
  1025 => (x"47",x"4f",x"52",x"50"),
  1026 => (x"2c",x"4d",x"41",x"52"),
  1027 => (x"4d",x"4f",x"53",x"20"),
  1028 => (x"54",x"53",x"20",x"45"),
  1029 => (x"47",x"4e",x"49",x"52"),
  1030 => (x"52",x"48",x"44",x"00"),
  1031 => (x"4f",x"54",x"53",x"59"),
  1032 => (x"50",x"20",x"45",x"4e"),
  1033 => (x"52",x"47",x"4f",x"52"),
  1034 => (x"20",x"2c",x"4d",x"41"),
  1035 => (x"54",x"53",x"27",x"31"),
  1036 => (x"52",x"54",x"53",x"20"),
  1037 => (x"00",x"47",x"4e",x"49"),
  1038 => (x"68",x"44",x"00",x"0a"),
  1039 => (x"74",x"73",x"79",x"72"),
  1040 => (x"20",x"65",x"6e",x"6f"),
  1041 => (x"63",x"6e",x"65",x"42"),
  1042 => (x"72",x"61",x"6d",x"68"),
  1043 => (x"56",x"20",x"2c",x"6b"),
  1044 => (x"69",x"73",x"72",x"65"),
  1045 => (x"32",x"20",x"6e",x"6f"),
  1046 => (x"28",x"20",x"31",x"2e"),
  1047 => (x"67",x"6e",x"61",x"4c"),
  1048 => (x"65",x"67",x"61",x"75"),
  1049 => (x"29",x"43",x"20",x"3a"),
  1050 => (x"00",x"0a",x"00",x"0a"),
  1051 => (x"63",x"65",x"78",x"45"),
  1052 => (x"6f",x"69",x"74",x"75"),
  1053 => (x"74",x"73",x"20",x"6e"),
  1054 => (x"73",x"74",x"72",x"61"),
  1055 => (x"64",x"25",x"20",x"2c"),
  1056 => (x"6e",x"75",x"72",x"20"),
  1057 => (x"68",x"74",x"20",x"73"),
  1058 => (x"67",x"75",x"6f",x"72"),
  1059 => (x"68",x"44",x"20",x"68"),
  1060 => (x"74",x"73",x"79",x"72"),
  1061 => (x"0a",x"65",x"6e",x"6f"),
  1062 => (x"65",x"78",x"45",x"00"),
  1063 => (x"69",x"74",x"75",x"63"),
  1064 => (x"65",x"20",x"6e",x"6f"),
  1065 => (x"0a",x"73",x"64",x"6e"),
  1066 => (x"46",x"00",x"0a",x"00"),
  1067 => (x"6c",x"61",x"6e",x"69"),
  1068 => (x"6c",x"61",x"76",x"20"),
  1069 => (x"20",x"73",x"65",x"75"),
  1070 => (x"74",x"20",x"66",x"6f"),
  1071 => (x"76",x"20",x"65",x"68"),
  1072 => (x"61",x"69",x"72",x"61"),
  1073 => (x"73",x"65",x"6c",x"62"),
  1074 => (x"65",x"73",x"75",x"20"),
  1075 => (x"6e",x"69",x"20",x"64"),
  1076 => (x"65",x"68",x"74",x"20"),
  1077 => (x"6e",x"65",x"62",x"20"),
  1078 => (x"61",x"6d",x"68",x"63"),
  1079 => (x"0a",x"3a",x"6b",x"72"),
  1080 => (x"49",x"00",x"0a",x"00"),
  1081 => (x"47",x"5f",x"74",x"6e"),
  1082 => (x"3a",x"62",x"6f",x"6c"),
  1083 => (x"20",x"20",x"20",x"20"),
  1084 => (x"20",x"20",x"20",x"20"),
  1085 => (x"20",x"20",x"20",x"20"),
  1086 => (x"00",x"0a",x"64",x"25"),
  1087 => (x"20",x"20",x"20",x"20"),
  1088 => (x"20",x"20",x"20",x"20"),
  1089 => (x"75",x"6f",x"68",x"73"),
  1090 => (x"62",x"20",x"64",x"6c"),
  1091 => (x"20",x"20",x"3a",x"65"),
  1092 => (x"0a",x"64",x"25",x"20"),
  1093 => (x"6f",x"6f",x"42",x"00"),
  1094 => (x"6c",x"47",x"5f",x"6c"),
  1095 => (x"20",x"3a",x"62",x"6f"),
  1096 => (x"20",x"20",x"20",x"20"),
  1097 => (x"20",x"20",x"20",x"20"),
  1098 => (x"64",x"25",x"20",x"20"),
  1099 => (x"20",x"20",x"00",x"0a"),
  1100 => (x"20",x"20",x"20",x"20"),
  1101 => (x"68",x"73",x"20",x"20"),
  1102 => (x"64",x"6c",x"75",x"6f"),
  1103 => (x"3a",x"65",x"62",x"20"),
  1104 => (x"25",x"20",x"20",x"20"),
  1105 => (x"43",x"00",x"0a",x"64"),
  1106 => (x"5f",x"31",x"5f",x"68"),
  1107 => (x"62",x"6f",x"6c",x"47"),
  1108 => (x"20",x"20",x"20",x"3a"),
  1109 => (x"20",x"20",x"20",x"20"),
  1110 => (x"20",x"20",x"20",x"20"),
  1111 => (x"00",x"0a",x"63",x"25"),
  1112 => (x"20",x"20",x"20",x"20"),
  1113 => (x"20",x"20",x"20",x"20"),
  1114 => (x"75",x"6f",x"68",x"73"),
  1115 => (x"62",x"20",x"64",x"6c"),
  1116 => (x"20",x"20",x"3a",x"65"),
  1117 => (x"0a",x"63",x"25",x"20"),
  1118 => (x"5f",x"68",x"43",x"00"),
  1119 => (x"6c",x"47",x"5f",x"32"),
  1120 => (x"20",x"3a",x"62",x"6f"),
  1121 => (x"20",x"20",x"20",x"20"),
  1122 => (x"20",x"20",x"20",x"20"),
  1123 => (x"63",x"25",x"20",x"20"),
  1124 => (x"20",x"20",x"00",x"0a"),
  1125 => (x"20",x"20",x"20",x"20"),
  1126 => (x"68",x"73",x"20",x"20"),
  1127 => (x"64",x"6c",x"75",x"6f"),
  1128 => (x"3a",x"65",x"62",x"20"),
  1129 => (x"25",x"20",x"20",x"20"),
  1130 => (x"41",x"00",x"0a",x"63"),
  1131 => (x"31",x"5f",x"72",x"72"),
  1132 => (x"6f",x"6c",x"47",x"5f"),
  1133 => (x"5d",x"38",x"5b",x"62"),
  1134 => (x"20",x"20",x"20",x"3a"),
  1135 => (x"20",x"20",x"20",x"20"),
  1136 => (x"00",x"0a",x"64",x"25"),
  1137 => (x"20",x"20",x"20",x"20"),
  1138 => (x"20",x"20",x"20",x"20"),
  1139 => (x"75",x"6f",x"68",x"73"),
  1140 => (x"62",x"20",x"64",x"6c"),
  1141 => (x"20",x"20",x"3a",x"65"),
  1142 => (x"0a",x"64",x"25",x"20"),
  1143 => (x"72",x"72",x"41",x"00"),
  1144 => (x"47",x"5f",x"32",x"5f"),
  1145 => (x"5b",x"62",x"6f",x"6c"),
  1146 => (x"37",x"5b",x"5d",x"38"),
  1147 => (x"20",x"20",x"3a",x"5d"),
  1148 => (x"64",x"25",x"20",x"20"),
  1149 => (x"20",x"20",x"00",x"0a"),
  1150 => (x"20",x"20",x"20",x"20"),
  1151 => (x"68",x"73",x"20",x"20"),
  1152 => (x"64",x"6c",x"75",x"6f"),
  1153 => (x"3a",x"65",x"62",x"20"),
  1154 => (x"4e",x"20",x"20",x"20"),
  1155 => (x"65",x"62",x"6d",x"75"),
  1156 => (x"66",x"4f",x"5f",x"72"),
  1157 => (x"6e",x"75",x"52",x"5f"),
  1158 => (x"20",x"2b",x"20",x"73"),
  1159 => (x"00",x"0a",x"30",x"31"),
  1160 => (x"5f",x"72",x"74",x"50"),
  1161 => (x"62",x"6f",x"6c",x"47"),
  1162 => (x"00",x"0a",x"3e",x"2d"),
  1163 => (x"74",x"50",x"20",x"20"),
  1164 => (x"6f",x"43",x"5f",x"72"),
  1165 => (x"20",x"3a",x"70",x"6d"),
  1166 => (x"20",x"20",x"20",x"20"),
  1167 => (x"20",x"20",x"20",x"20"),
  1168 => (x"0a",x"64",x"25",x"20"),
  1169 => (x"20",x"20",x"20",x"00"),
  1170 => (x"20",x"20",x"20",x"20"),
  1171 => (x"6f",x"68",x"73",x"20"),
  1172 => (x"20",x"64",x"6c",x"75"),
  1173 => (x"20",x"3a",x"65",x"62"),
  1174 => (x"69",x"28",x"20",x"20"),
  1175 => (x"65",x"6c",x"70",x"6d"),
  1176 => (x"74",x"6e",x"65",x"6d"),
  1177 => (x"6f",x"69",x"74",x"61"),
  1178 => (x"65",x"64",x"2d",x"6e"),
  1179 => (x"64",x"6e",x"65",x"70"),
  1180 => (x"29",x"74",x"6e",x"65"),
  1181 => (x"20",x"20",x"00",x"0a"),
  1182 => (x"63",x"73",x"69",x"44"),
  1183 => (x"20",x"20",x"3a",x"72"),
  1184 => (x"20",x"20",x"20",x"20"),
  1185 => (x"20",x"20",x"20",x"20"),
  1186 => (x"25",x"20",x"20",x"20"),
  1187 => (x"20",x"00",x"0a",x"64"),
  1188 => (x"20",x"20",x"20",x"20"),
  1189 => (x"73",x"20",x"20",x"20"),
  1190 => (x"6c",x"75",x"6f",x"68"),
  1191 => (x"65",x"62",x"20",x"64"),
  1192 => (x"20",x"20",x"20",x"3a"),
  1193 => (x"00",x"0a",x"64",x"25"),
  1194 => (x"6e",x"45",x"20",x"20"),
  1195 => (x"43",x"5f",x"6d",x"75"),
  1196 => (x"3a",x"70",x"6d",x"6f"),
  1197 => (x"20",x"20",x"20",x"20"),
  1198 => (x"20",x"20",x"20",x"20"),
  1199 => (x"0a",x"64",x"25",x"20"),
  1200 => (x"20",x"20",x"20",x"00"),
  1201 => (x"20",x"20",x"20",x"20"),
  1202 => (x"6f",x"68",x"73",x"20"),
  1203 => (x"20",x"64",x"6c",x"75"),
  1204 => (x"20",x"3a",x"65",x"62"),
  1205 => (x"64",x"25",x"20",x"20"),
  1206 => (x"20",x"20",x"00",x"0a"),
  1207 => (x"5f",x"74",x"6e",x"49"),
  1208 => (x"70",x"6d",x"6f",x"43"),
  1209 => (x"20",x"20",x"20",x"3a"),
  1210 => (x"20",x"20",x"20",x"20"),
  1211 => (x"25",x"20",x"20",x"20"),
  1212 => (x"20",x"00",x"0a",x"64"),
  1213 => (x"20",x"20",x"20",x"20"),
  1214 => (x"73",x"20",x"20",x"20"),
  1215 => (x"6c",x"75",x"6f",x"68"),
  1216 => (x"65",x"62",x"20",x"64"),
  1217 => (x"20",x"20",x"20",x"3a"),
  1218 => (x"00",x"0a",x"64",x"25"),
  1219 => (x"74",x"53",x"20",x"20"),
  1220 => (x"6f",x"43",x"5f",x"72"),
  1221 => (x"20",x"3a",x"70",x"6d"),
  1222 => (x"20",x"20",x"20",x"20"),
  1223 => (x"20",x"20",x"20",x"20"),
  1224 => (x"0a",x"73",x"25",x"20"),
  1225 => (x"20",x"20",x"20",x"00"),
  1226 => (x"20",x"20",x"20",x"20"),
  1227 => (x"6f",x"68",x"73",x"20"),
  1228 => (x"20",x"64",x"6c",x"75"),
  1229 => (x"20",x"3a",x"65",x"62"),
  1230 => (x"48",x"44",x"20",x"20"),
  1231 => (x"54",x"53",x"59",x"52"),
  1232 => (x"20",x"45",x"4e",x"4f"),
  1233 => (x"47",x"4f",x"52",x"50"),
  1234 => (x"2c",x"4d",x"41",x"52"),
  1235 => (x"4d",x"4f",x"53",x"20"),
  1236 => (x"54",x"53",x"20",x"45"),
  1237 => (x"47",x"4e",x"49",x"52"),
  1238 => (x"65",x"4e",x"00",x"0a"),
  1239 => (x"50",x"5f",x"74",x"78"),
  1240 => (x"47",x"5f",x"72",x"74"),
  1241 => (x"2d",x"62",x"6f",x"6c"),
  1242 => (x"20",x"00",x"0a",x"3e"),
  1243 => (x"72",x"74",x"50",x"20"),
  1244 => (x"6d",x"6f",x"43",x"5f"),
  1245 => (x"20",x"20",x"3a",x"70"),
  1246 => (x"20",x"20",x"20",x"20"),
  1247 => (x"20",x"20",x"20",x"20"),
  1248 => (x"00",x"0a",x"64",x"25"),
  1249 => (x"20",x"20",x"20",x"20"),
  1250 => (x"20",x"20",x"20",x"20"),
  1251 => (x"75",x"6f",x"68",x"73"),
  1252 => (x"62",x"20",x"64",x"6c"),
  1253 => (x"20",x"20",x"3a",x"65"),
  1254 => (x"6d",x"69",x"28",x"20"),
  1255 => (x"6d",x"65",x"6c",x"70"),
  1256 => (x"61",x"74",x"6e",x"65"),
  1257 => (x"6e",x"6f",x"69",x"74"),
  1258 => (x"70",x"65",x"64",x"2d"),
  1259 => (x"65",x"64",x"6e",x"65"),
  1260 => (x"2c",x"29",x"74",x"6e"),
  1261 => (x"6d",x"61",x"73",x"20"),
  1262 => (x"73",x"61",x"20",x"65"),
  1263 => (x"6f",x"62",x"61",x"20"),
  1264 => (x"00",x"0a",x"65",x"76"),
  1265 => (x"69",x"44",x"20",x"20"),
  1266 => (x"3a",x"72",x"63",x"73"),
  1267 => (x"20",x"20",x"20",x"20"),
  1268 => (x"20",x"20",x"20",x"20"),
  1269 => (x"20",x"20",x"20",x"20"),
  1270 => (x"0a",x"64",x"25",x"20"),
  1271 => (x"20",x"20",x"20",x"00"),
  1272 => (x"20",x"20",x"20",x"20"),
  1273 => (x"6f",x"68",x"73",x"20"),
  1274 => (x"20",x"64",x"6c",x"75"),
  1275 => (x"20",x"3a",x"65",x"62"),
  1276 => (x"64",x"25",x"20",x"20"),
  1277 => (x"20",x"20",x"00",x"0a"),
  1278 => (x"6d",x"75",x"6e",x"45"),
  1279 => (x"6d",x"6f",x"43",x"5f"),
  1280 => (x"20",x"20",x"3a",x"70"),
  1281 => (x"20",x"20",x"20",x"20"),
  1282 => (x"25",x"20",x"20",x"20"),
  1283 => (x"20",x"00",x"0a",x"64"),
  1284 => (x"20",x"20",x"20",x"20"),
  1285 => (x"73",x"20",x"20",x"20"),
  1286 => (x"6c",x"75",x"6f",x"68"),
  1287 => (x"65",x"62",x"20",x"64"),
  1288 => (x"20",x"20",x"20",x"3a"),
  1289 => (x"00",x"0a",x"64",x"25"),
  1290 => (x"6e",x"49",x"20",x"20"),
  1291 => (x"6f",x"43",x"5f",x"74"),
  1292 => (x"20",x"3a",x"70",x"6d"),
  1293 => (x"20",x"20",x"20",x"20"),
  1294 => (x"20",x"20",x"20",x"20"),
  1295 => (x"0a",x"64",x"25",x"20"),
  1296 => (x"20",x"20",x"20",x"00"),
  1297 => (x"20",x"20",x"20",x"20"),
  1298 => (x"6f",x"68",x"73",x"20"),
  1299 => (x"20",x"64",x"6c",x"75"),
  1300 => (x"20",x"3a",x"65",x"62"),
  1301 => (x"64",x"25",x"20",x"20"),
  1302 => (x"20",x"20",x"00",x"0a"),
  1303 => (x"5f",x"72",x"74",x"53"),
  1304 => (x"70",x"6d",x"6f",x"43"),
  1305 => (x"20",x"20",x"20",x"3a"),
  1306 => (x"20",x"20",x"20",x"20"),
  1307 => (x"25",x"20",x"20",x"20"),
  1308 => (x"20",x"00",x"0a",x"73"),
  1309 => (x"20",x"20",x"20",x"20"),
  1310 => (x"73",x"20",x"20",x"20"),
  1311 => (x"6c",x"75",x"6f",x"68"),
  1312 => (x"65",x"62",x"20",x"64"),
  1313 => (x"20",x"20",x"20",x"3a"),
  1314 => (x"59",x"52",x"48",x"44"),
  1315 => (x"4e",x"4f",x"54",x"53"),
  1316 => (x"52",x"50",x"20",x"45"),
  1317 => (x"41",x"52",x"47",x"4f"),
  1318 => (x"53",x"20",x"2c",x"4d"),
  1319 => (x"20",x"45",x"4d",x"4f"),
  1320 => (x"49",x"52",x"54",x"53"),
  1321 => (x"00",x"0a",x"47",x"4e"),
  1322 => (x"5f",x"74",x"6e",x"49"),
  1323 => (x"6f",x"4c",x"5f",x"31"),
  1324 => (x"20",x"20",x"3a",x"63"),
  1325 => (x"20",x"20",x"20",x"20"),
  1326 => (x"20",x"20",x"20",x"20"),
  1327 => (x"0a",x"64",x"25",x"20"),
  1328 => (x"20",x"20",x"20",x"00"),
  1329 => (x"20",x"20",x"20",x"20"),
  1330 => (x"6f",x"68",x"73",x"20"),
  1331 => (x"20",x"64",x"6c",x"75"),
  1332 => (x"20",x"3a",x"65",x"62"),
  1333 => (x"64",x"25",x"20",x"20"),
  1334 => (x"6e",x"49",x"00",x"0a"),
  1335 => (x"5f",x"32",x"5f",x"74"),
  1336 => (x"3a",x"63",x"6f",x"4c"),
  1337 => (x"20",x"20",x"20",x"20"),
  1338 => (x"20",x"20",x"20",x"20"),
  1339 => (x"25",x"20",x"20",x"20"),
  1340 => (x"20",x"00",x"0a",x"64"),
  1341 => (x"20",x"20",x"20",x"20"),
  1342 => (x"73",x"20",x"20",x"20"),
  1343 => (x"6c",x"75",x"6f",x"68"),
  1344 => (x"65",x"62",x"20",x"64"),
  1345 => (x"20",x"20",x"20",x"3a"),
  1346 => (x"00",x"0a",x"64",x"25"),
  1347 => (x"5f",x"74",x"6e",x"49"),
  1348 => (x"6f",x"4c",x"5f",x"33"),
  1349 => (x"20",x"20",x"3a",x"63"),
  1350 => (x"20",x"20",x"20",x"20"),
  1351 => (x"20",x"20",x"20",x"20"),
  1352 => (x"0a",x"64",x"25",x"20"),
  1353 => (x"20",x"20",x"20",x"00"),
  1354 => (x"20",x"20",x"20",x"20"),
  1355 => (x"6f",x"68",x"73",x"20"),
  1356 => (x"20",x"64",x"6c",x"75"),
  1357 => (x"20",x"3a",x"65",x"62"),
  1358 => (x"64",x"25",x"20",x"20"),
  1359 => (x"6e",x"45",x"00",x"0a"),
  1360 => (x"4c",x"5f",x"6d",x"75"),
  1361 => (x"20",x"3a",x"63",x"6f"),
  1362 => (x"20",x"20",x"20",x"20"),
  1363 => (x"20",x"20",x"20",x"20"),
  1364 => (x"25",x"20",x"20",x"20"),
  1365 => (x"20",x"00",x"0a",x"64"),
  1366 => (x"20",x"20",x"20",x"20"),
  1367 => (x"73",x"20",x"20",x"20"),
  1368 => (x"6c",x"75",x"6f",x"68"),
  1369 => (x"65",x"62",x"20",x"64"),
  1370 => (x"20",x"20",x"20",x"3a"),
  1371 => (x"00",x"0a",x"64",x"25"),
  1372 => (x"5f",x"72",x"74",x"53"),
  1373 => (x"6f",x"4c",x"5f",x"31"),
  1374 => (x"20",x"20",x"3a",x"63"),
  1375 => (x"20",x"20",x"20",x"20"),
  1376 => (x"20",x"20",x"20",x"20"),
  1377 => (x"0a",x"73",x"25",x"20"),
  1378 => (x"20",x"20",x"20",x"00"),
  1379 => (x"20",x"20",x"20",x"20"),
  1380 => (x"6f",x"68",x"73",x"20"),
  1381 => (x"20",x"64",x"6c",x"75"),
  1382 => (x"20",x"3a",x"65",x"62"),
  1383 => (x"48",x"44",x"20",x"20"),
  1384 => (x"54",x"53",x"59",x"52"),
  1385 => (x"20",x"45",x"4e",x"4f"),
  1386 => (x"47",x"4f",x"52",x"50"),
  1387 => (x"2c",x"4d",x"41",x"52"),
  1388 => (x"53",x"27",x"31",x"20"),
  1389 => (x"54",x"53",x"20",x"54"),
  1390 => (x"47",x"4e",x"49",x"52"),
  1391 => (x"74",x"53",x"00",x"0a"),
  1392 => (x"5f",x"32",x"5f",x"72"),
  1393 => (x"3a",x"63",x"6f",x"4c"),
  1394 => (x"20",x"20",x"20",x"20"),
  1395 => (x"20",x"20",x"20",x"20"),
  1396 => (x"25",x"20",x"20",x"20"),
  1397 => (x"20",x"00",x"0a",x"73"),
  1398 => (x"20",x"20",x"20",x"20"),
  1399 => (x"73",x"20",x"20",x"20"),
  1400 => (x"6c",x"75",x"6f",x"68"),
  1401 => (x"65",x"62",x"20",x"64"),
  1402 => (x"20",x"20",x"20",x"3a"),
  1403 => (x"59",x"52",x"48",x"44"),
  1404 => (x"4e",x"4f",x"54",x"53"),
  1405 => (x"52",x"50",x"20",x"45"),
  1406 => (x"41",x"52",x"47",x"4f"),
  1407 => (x"32",x"20",x"2c",x"4d"),
  1408 => (x"20",x"44",x"4e",x"27"),
  1409 => (x"49",x"52",x"54",x"53"),
  1410 => (x"00",x"0a",x"47",x"4e"),
  1411 => (x"73",x"55",x"00",x"0a"),
  1412 => (x"74",x"20",x"72",x"65"),
  1413 => (x"3a",x"65",x"6d",x"69"),
  1414 => (x"0a",x"64",x"25",x"20"),
  1415 => (x"00",x"00",x"00",x"00"),
  1416 => (x"d0",x"90",x"00",x"00"),
  1417 => (x"d0",x"90",x"00",x"03"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Xilinx XST attributes
	attribute ram_style: string;
	attribute ram_style of ram: signal is "no_rw_check";

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(from_soc.memAAddr(maxAddrBitBRAM downto 2)));

	-- Reorganize the read data from the RAM to match the output
	unpack: for i in 0 to BYTES - 1 generate    
		data_out1(BYTE_WIDTH*(i+1) - 1 downto BYTE_WIDTH*i) <= q1_local((BYTES-1)-i);
	end generate unpack;
        
	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we1 = '1') then
				-- edit this code if using other than four bytes per word
				if(be1(3) = '1') then
					ram(addr1)(3) <= data_in1(7 downto 0);
				end if;
				if be1(2) = '1' then
					ram(addr1)(2) <= data_in1(15 downto 8);
				end if;
				if be1(1) = '1' then
					ram(addr1)(1) <= data_in1(23 downto 16);
				end if;
				if be1(0) = '1' then
					ram(addr1)(0) <= data_in1(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;
